/*Copyright 2020-2021 T-Head Semiconductor Co., Ltd.

Licensed under the Apache License, Version 2.0 (the "License");
you may not use this file except in compliance with the License.
You may obtain a copy of the License at

    http://www.apache.org/licenses/LICENSE-2.0

Unless required by applicable law or agreed to in writing, software
distributed under the License is distributed on an "AS IS" BASIS,
WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
See the License for the specific language governing permissions and
limitations under the License.
*/

// &ModuleBeg; @22
module aq_spsram_128x8(
  A,
  CEN,
  CLK,
  D,
  GWEN,
  Q,
  WEN
);

// &Ports; @23
input   [6:0]  A;   
input          CEN; 
input          CLK; 
input   [7:0]  D;   
input          GWEN; 
input   [7:0]  WEN; 
output  [7:0]  Q;   

// &Regs; @24

// &Wires; @25
wire    [6:0]  A;   
wire           CEN; 
wire           CLK; 
wire    [7:0]  D;   
wire           GWEN; 
wire    [7:0]  Q;   
wire    [7:0]  WEN; 


//**********************************************************
//                  Parameter Definition
//**********************************************************
parameter ADDR_WIDTH = 7;
parameter DATA_WIDTH = 8;
parameter WE_WIDTH   = 8;

//  //********************************************************
//  //*                        FPGA memory                   *
//  //********************************************************
//   &Instance("aq_f_spsram_128x8"); @43
aq_f_spsram_128x8  x_aq_f_spsram_128x8 (
  .A    (A   ),
  .CEN  (CEN ),
  .CLK  (CLK ),
  .D    (D   ),
  .GWEN (GWEN),
  .Q    (Q   ),
  .WEN  (WEN )
);

endmodule



